
int num_errors = 0;
